--------------------
-- 4096*16 Memory --
--------------------
ENTITY memory IS
    PORT
    (
        i : IN bit_vector(15 DOWNTO 0);
        a : IN bit_vector(11 DOWNTO 0);
        rm,wm,clock : IN bit;
        o : OUT bit_vector(15 DOWNTO 0)
    );
END memory;

ARCHITECTURE memory_arch OF memory IS
    FUNCTION convert (x : bit_vector) RETURN integer IS
    VARIABLE sum : integer:=0;
    VARIABLE j : integer;
    BEGIN
        FOR j IN x'RANGE LOOP
            IF x(j)='1' THEN
                sum := sum + 2**j;
            END IF;
        END LOOP;
        RETURN sum;
    END convert;
    TYPE ram_type IS ARRAY (4095 DOWNTO 0) OF bit_vector(15 DOWNTO 0);
    SIGNAL ram : ram_type:=
        (
                 0 => "0111000000000100",
                 1 => "0100000011001000",
                 2 => "0100000000000011",
                 3 => "0010000001100100",
                 4 => "0111001000000000",
                 5 => "0111000000100000",
                 6 => "0101000000010011",
                 7 => "0111000000000001",
                20 => "1001000001100101",
                21 => "0111000000010000",
                22 => "0100000000011010",
                23 => "0111000010000000",
                24 => "0000000001101010",
                25 => "0100000000100000",
                26 => "0111000010000000",
                27 => "0111000000000010",
                28 => "0100000000100000",
                29 => "0111001000000000",
                30 => "0000000001101010",
                31 => "0111001000000000",
                32 => "0110000001100111",
                33 => "0100000000010101",
                34 => "1111000100000000",
                35 => "0100000000100010",
                36 => "1111010000000000",
                37 => "1011000001101000",
                38 => "1001000001100101",
                39 => "1111000010000000",
                40 => "1100000000010011",
               100 => "0000000010100010",
               101 => "0000000001100110",
               102 => "0000000000000010",
               103 => "1111111111111100",
               104 => "0000000001101001",
               106 => "0111111111111111",
               200 => "1111000100000000",
               201 => "0100000011001011",
               202 => "1111010000000000",
               203 => "1111000010000000",
               204 => "1100000000000000",
            OTHERS => "0000000000000000"
        );
    BEGIN
        PROCESS(rm,wm,a,i,clock)
            BEGIN
                IF (clock'event AND clock='1') THEN
                    IF wm='1' THEN
                        ram(convert(a)) <= i;
                    END IF;
                END IF;
                IF rm='1' THEN
                    o <= ram(convert(a));
                END IF;
                IF rm='0' AND wm='0' THEN
                    NULL;
                END IF;
            END PROCESS;
    END memory_arch;