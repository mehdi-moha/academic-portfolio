* H:\Lab-5\lab-5-3\lab-5-3.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 17:34:04 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-5-3.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-5-3.net"
.INC "lab-5-3.als"


.probe


.END
