* H:\Lab-1\lab-1-2\lab-1-2.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 17:25:54 2005



** Analysis setup **
.tran 1ms 6ms
.OP 
.STMLIB "lab-1-2.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-1-2.net"
.INC "lab-1-2.als"


.probe


.END
