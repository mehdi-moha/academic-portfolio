* H:\Lab-4\lab-4-1\lab-4-1.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 10:53:03 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-4-1.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-4-1.net"
.INC "lab-4-1.als"


.probe


.END
