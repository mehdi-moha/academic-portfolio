* H:\Lab-1\lab-1-5\lab-1-5-4081.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 18:01:19 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-1-5-4081.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-1-5-4081.net"
.INC "lab-1-5-4081.als"


.probe


.END
