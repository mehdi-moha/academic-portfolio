* H:\Lab-3\lab-3-5\lab-3-5.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 15:54:47 2005



** Analysis setup **
.tran 1ms 10ms
.OP 
.STMLIB "lab-3-5.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-3-5.net"
.INC "lab-3-5.als"


.probe


.END
