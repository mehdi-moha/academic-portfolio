* H:\Lab-4\lab-4-2\lab-4-2.sch

* Schematics Version 9.1 - Web Update 1
* Sun May 29 01:02:23 2005



** Analysis setup **
.tran 1ms 6ms
.OP 
.STMLIB "lab-4-2.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-4-2.net"
.INC "lab-4-2.als"


.probe


.END
