* H:\Lab-1\lab-1-1\lab-1-1.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 17:32:06 2005



** Analysis setup **
.tran 1ms 6ms
.OP 
.STMLIB "lab-1-1.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-1-1.net"
.INC "lab-1-1.als"


.probe


.END
