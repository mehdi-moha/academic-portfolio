* H:\Lab-2\Lab-2-1\nor\nor.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 15:23:55 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "nor.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "nor.net"
.INC "nor.als"


.probe


.END
