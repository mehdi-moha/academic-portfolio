* H:\Lab-4\lab-4-4\lab-4-4.sch

* Schematics Version 9.1 - Web Update 1
* Sun May 29 20:27:54 2005



** Analysis setup **
.tran 1ms 6ms
.OP 


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-4-4.net"
.INC "lab-4-4.als"


.probe


.END
