* H:\Lab-5\lab-5-1\lab-5-1.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 21:24:36 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-5-1.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-5-1.net"
.INC "lab-5-1.als"


.probe


.END
