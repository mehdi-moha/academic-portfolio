* H:\Lab-3\lab-3-1\lab-3-1.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 08:02:39 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-3-1.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-3-1.net"
.INC "lab-3-1.als"


.probe


.END
