* H:\Lab-2\Lab-2-1\or\or.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 13:09:28 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "or.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "or.net"
.INC "or.als"


.probe


.END
