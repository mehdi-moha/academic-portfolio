* H:\Lab-1\lab-1-4-t4\lab-1-4-t4.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 17:41:06 2005



** Analysis setup **
.tran 1ms 10ms
.OP 
.STMLIB "lab-1-4-t4.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-1-4-t4.net"
.INC "lab-1-4-t4.als"


.probe


.END
