* H:\Lab-1\lab-1-4\lab-1-4.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 28 17:31:13 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-1-4.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-1-4.net"
.INC "lab-1-4.als"


.probe


.END
