* H:\Lab-2\Q-2\nand-xor\xor.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 15:44:16 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "xor.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "xor.net"
.INC "xor.als"


.probe


.END
