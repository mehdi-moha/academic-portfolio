* H:\Lab-7\lab-7-1\lab-7-1.sch

* Schematics Version 9.1 - Web Update 1
* Mon May 30 17:08:21 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "lab-7-1.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-7-1.net"
.INC "lab-7-1.als"


.probe


.END
