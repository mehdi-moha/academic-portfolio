* H:\Lab-2\Lab-2-3\nand\nand.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 15:23:00 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "nand.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "nand.net"
.INC "nand.als"


.probe


.END
