* H:\Lab-4\lab-4-2-6bit\lab-4-2-6bit.sch

* Schematics Version 9.1 - Web Update 1
* Sun May 29 19:35:33 2005



** Analysis setup **
.tran 1ms 6ms
.OP 
.STMLIB "lab-4-2-6bit.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "lab-4-2-6bit.net"
.INC "lab-4-2-6bit.als"


.probe


.END
