* H:\Lab-2\Lab-2-1\not\not.sch

* Schematics Version 9.1 - Web Update 1
* Fri May 27 15:24:39 2005



** Analysis setup **
.tran 1ms 8ms
.OP 
.STMLIB "not.stl"


* From [PSPICE NETLIST] section of pspice91.ini:
.lib "nom.lib"

.INC "not.net"
.INC "not.als"


.probe


.END
